library IEEE;
use IEEE.std_logic_1164.ALL;

entity rowselect1 is
   port(a :in    std_logic_vector(5 downto 0);
        c1:out   std_logic);
end rowselect1;