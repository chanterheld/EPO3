architecture behav of rng is 

begin


end behav;
