library ieee;
use ieee.std_logic_1164.all;

entity seg_10 is
	port(	a	: in	std_logic;
		b	: in	std_logic;
		c	: in	std_logic;
		d	: in	std_logic;
		state 	: out	std_logic
	);
end seg_10;